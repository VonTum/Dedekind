`timescale 1ns / 1ps

module testPermuteCheck720();

reg clk = 0;
initial forever #1 clk = !clk;



endmodule
